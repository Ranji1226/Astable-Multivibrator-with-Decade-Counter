* /home/sranjith102001/Desktop/ranji_esim/ranji_decade_counter/ranji_decade_counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 09 Mar 2022 06:08:30 PM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_R1-Pad1_ Net-_C1-Pad2_ 510		
R2  Net-_R1-Pad1_ Net-_C2-Pad2_ 10k		
R3  Net-_R1-Pad1_ Net-_C1-Pad1_ 10k		
R4  Net-_R1-Pad1_ Out 510		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 100u		
C2  Out Net-_C2-Pad2_ 100u		
Q2  Out Net-_C1-Pad1_ GND eSim_NPN		
Q1  Net-_C1-Pad2_ Net-_C2-Pad2_ GND eSim_NPN		
U3  Net-_U3-Pad1_ Out Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
U4  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ O1 o2 o3 o4 dac_bridge_4		
v1  Net-_R1-Pad1_ GND DC		
v2  GND Net-_U3-Pad1_ pulse		
U1  ? plot_v1		
U5  O1 plot_v1		
U6  o2 plot_v1		
U7  o3 plot_v1		
U8  o4 plot_v1		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ ranji_decadecounter		

.end
